
module caliptra_ss_package_top (
    input wire core_clk,
    input wire rst_l,
    input wire porst_l,
    /*
    // Caliptra AXI Interface
    input  wire [31:0] S_AXI_CALIPTRA_AWADDR,
    input  wire [1:0] S_AXI_CALIPTRA_AWBURST,
    input  wire [2:0] S_AXI_CALIPTRA_AWSIZE,
    input  wire [7:0] S_AXI_CALIPTRA_AWLEN,
    input  wire [31:0] S_AXI_CALIPTRA_AWUSER,
    input  wire [15:0] S_AXI_CALIPTRA_AWID,
    input  wire S_AXI_CALIPTRA_AWLOCK,
    input  wire S_AXI_CALIPTRA_AWVALID,
    output wire S_AXI_CALIPTRA_AWREADY,
    // W
    input  wire [31:0] S_AXI_CALIPTRA_WDATA,
    input  wire [3:0] S_AXI_CALIPTRA_WSTRB,
    input  wire S_AXI_CALIPTRA_WVALID,
    output wire S_AXI_CALIPTRA_WREADY,
    input  wire S_AXI_CALIPTRA_WLAST,
    // B
    output wire [1:0] S_AXI_CALIPTRA_BRESP,
    output reg  [15:0] S_AXI_CALIPTRA_BID,
    output wire S_AXI_CALIPTRA_BVALID,
    input  wire S_AXI_CALIPTRA_BREADY,
    // AR
    input  wire [31:0] S_AXI_CALIPTRA_ARADDR,
    input  wire [1:0] S_AXI_CALIPTRA_ARBURST,
    input  wire [2:0] S_AXI_CALIPTRA_ARSIZE,
    input  wire [7:0] S_AXI_CALIPTRA_ARLEN,
    input  wire [31:0] S_AXI_CALIPTRA_ARUSER,
    input  wire [15:0] S_AXI_CALIPTRA_ARID,
    input  wire S_AXI_CALIPTRA_ARLOCK,
    input  wire S_AXI_CALIPTRA_ARVALID,
    output wire S_AXI_CALIPTRA_ARREADY,
    // R
    output wire [31:0] S_AXI_CALIPTRA_RDATA,
    output wire [3:0] S_AXI_CALIPTRA_RRESP,
    output reg  [15:0] S_AXI_CALIPTRA_RID,
    output wire S_AXI_CALIPTRA_RLAST,
    output wire S_AXI_CALIPTRA_RVALID,
    input  wire S_AXI_CALIPTRA_RREADY,
*/
    //-------------------------- LSU AXI signals--------------------------
    // AXI Write Channels
    output wire                      M_AXI_MCU_LSU_AWVALID,
    input  wire                      M_AXI_MCU_LSU_AWREADY,
    output wire [3-1:0]              M_AXI_MCU_LSU_AWID,
    output wire [              31:0] M_AXI_MCU_LSU_AWADDR,
    output wire [               3:0] M_AXI_MCU_LSU_AWREGION,
    output wire [               7:0] M_AXI_MCU_LSU_AWLEN,
    output wire [               2:0] M_AXI_MCU_LSU_AWSIZE,
    output wire [               1:0] M_AXI_MCU_LSU_AWBURST,
    output wire                      M_AXI_MCU_LSU_AWLOCK,
    output wire [               3:0] M_AXI_MCU_LSU_AWCACHE,
    output wire [               2:0] M_AXI_MCU_LSU_AWPROT,
    output wire [               3:0] M_AXI_MCU_LSU_AWQOS,

    output wire                      M_AXI_MCU_LSU_WVALID,
    input  wire                      M_AXI_MCU_LSU_WREADY,
    output wire [63:0]               M_AXI_MCU_LSU_WDATA,
    output wire [ 7:0]               M_AXI_MCU_LSU_WSTRB,
    output wire                      M_AXI_MCU_LSU_WLAST,

    input  wire                      M_AXI_MCU_LSU_BVALID,
    output wire                      M_AXI_MCU_LSU_BREADY,
    input  wire [               1:0] M_AXI_MCU_LSU_BRESP,
    input  wire [3-1:0]              M_AXI_MCU_LSU_BID,

    // AXI Read Channels
    output wire                      M_AXI_MCU_LSU_ARVALID,
    input  wire                      M_AXI_MCU_LSU_ARREADY,
    output wire [3-1:0]              M_AXI_MCU_LSU_ARID,
    output wire [              31:0] M_AXI_MCU_LSU_ARADDR,
    output wire [               3:0] M_AXI_MCU_LSU_ARREGION,
    output wire [               7:0] M_AXI_MCU_LSU_ARLEN,
    output wire [               2:0] M_AXI_MCU_LSU_ARSIZE,
    output wire [               1:0] M_AXI_MCU_LSU_ARBURST,
    output wire                      M_AXI_MCU_LSU_ARLOCK,
    output wire [               3:0] M_AXI_MCU_LSU_ARCACHE,
    output wire [               2:0] M_AXI_MCU_LSU_ARPROT,
    output wire [               3:0] M_AXI_MCU_LSU_ARQOS,

    input  wire                      M_AXI_MCU_LSU_RVALID,
    output wire                      M_AXI_MCU_LSU_RREADY,
    input  wire [3-1:0]              M_AXI_MCU_LSU_RID,
    input  wire [              63:0] M_AXI_MCU_LSU_RDATA,
    input  wire [               1:0] M_AXI_MCU_LSU_RRESP,
    input  wire                      M_AXI_MCU_LSU_RLAST,

    //-------------------------- IFU AXI signals--------------------------
    // AXI Write Channels
    output wire                      M_AXI_MCU_IFU_AWVALID,
    input  wire                      M_AXI_MCU_IFU_AWREADY,
    output wire [3-1:0]              M_AXI_MCU_IFU_AWID,
    output wire [              31:0] M_AXI_MCU_IFU_AWADDR,
    output wire [               3:0] M_AXI_MCU_IFU_AWREGION,
    output wire [               7:0] M_AXI_MCU_IFU_AWLEN,
    output wire [               2:0] M_AXI_MCU_IFU_AWSIZE,
    output wire [               1:0] M_AXI_MCU_IFU_AWBURST,
    output wire                      M_AXI_MCU_IFU_AWLOCK,
    output wire [               3:0] M_AXI_MCU_IFU_AWCACHE,
    output wire [               2:0] M_AXI_MCU_IFU_AWPROT,
    output wire [               3:0] M_AXI_MCU_IFU_AWQOS,

    output wire                      M_AXI_MCU_IFU_WVALID,
    input  wire                      M_AXI_MCU_IFU_WREADY,
    output wire [63:0]               M_AXI_MCU_IFU_WDATA,
    output wire [ 7:0]               M_AXI_MCU_IFU_WSTRB,
    output wire                      M_AXI_MCU_IFU_WLAST,

    input  wire                      M_AXI_MCU_IFU_BVALID,
    output wire                      M_AXI_MCU_IFU_BREADY,
    input  wire [               1:0] M_AXI_MCU_IFU_BRESP,
    input  wire [3-1:0]              M_AXI_MCU_IFU_BID,

    // AXI Read Channels
    output wire                      M_AXI_MCU_IFU_ARVALID,
    input  wire                      M_AXI_MCU_IFU_ARREADY,
    output wire [3-1:0]              M_AXI_MCU_IFU_ARID,
    output wire [              31:0] M_AXI_MCU_IFU_ARADDR,
    output wire [               3:0] M_AXI_MCU_IFU_ARREGION,
    output wire [               7:0] M_AXI_MCU_IFU_ARLEN,
    output wire [               2:0] M_AXI_MCU_IFU_ARSIZE,
    output wire [               1:0] M_AXI_MCU_IFU_ARBURST,
    output wire                      M_AXI_MCU_IFU_ARLOCK,
    output wire [               3:0] M_AXI_MCU_IFU_ARCACHE,
    output wire [               2:0] M_AXI_MCU_IFU_ARPROT,
    output wire [               3:0] M_AXI_MCU_IFU_ARQOS,

    input  wire                      M_AXI_MCU_IFU_RVALID,
    output wire                      M_AXI_MCU_IFU_RREADY,
    input  wire [3-1:0]              M_AXI_MCU_IFU_RID,
    input  wire [              63:0] M_AXI_MCU_IFU_RDATA,
    input  wire [               1:0] M_AXI_MCU_IFU_RRESP,
    input  wire                      M_AXI_MCU_IFU_RLAST,

    //-------------------------- SB AXI signals--------------------------
    // AXI Write Channels
    output wire                     sb_axi_awvalid,
    input  wire                     sb_axi_awready,
    output wire [1-1:0]             sb_axi_awid,
    output wire [             31:0] sb_axi_awaddr,
    output wire [              3:0] sb_axi_awregion,
    output wire [              7:0] sb_axi_awlen,
    output wire [              2:0] sb_axi_awsize,
    output wire [              1:0] sb_axi_awburst,
    output wire                     sb_axi_awlock,
    output wire [              3:0] sb_axi_awcache,
    output wire [              2:0] sb_axi_awprot,
    output wire [              3:0] sb_axi_awqos,

    output wire                     sb_axi_wvalid,
    input  wire                     sb_axi_wready,
    output wire [63:0]              sb_axi_wdata,
    output wire [ 7:0]              sb_axi_wstrb,
    output wire                     sb_axi_wlast,

    input  wire                     sb_axi_bvalid,
    output wire                     sb_axi_bready,
    input  wire [              1:0] sb_axi_bresp,
    input  wire [1-1:0]             sb_axi_bid,

    // AXI Read Channels
    output wire                     sb_axi_arvalid,
    input  wire                     sb_axi_arready,
    output wire [1-1:0]             sb_axi_arid,
    output wire [             31:0] sb_axi_araddr,
    output wire [              3:0] sb_axi_arregion,
    output wire [              7:0] sb_axi_arlen,
    output wire [              2:0] sb_axi_arsize,
    output wire [              1:0] sb_axi_arburst,
    output wire                     sb_axi_arlock,
    output wire [              3:0] sb_axi_arcache,
    output wire [              2:0] sb_axi_arprot,
    output wire [              3:0] sb_axi_arqos,

    input  wire                     sb_axi_rvalid,
    output wire                     sb_axi_rready,
    input  wire [1-1:0]             sb_axi_rid,
    input  wire [             63:0] sb_axi_rdata,
    input  wire [              1:0] sb_axi_rresp,
    input  wire                     sb_axi_rlast,

    //-------------------------- DMA AXI signals--------------------------
    // AXI Write Channels
    input  wire                      S_AXI_MCU_DMA_AWVALID,
    output wire                      S_AXI_MCU_DMA_AWREADY,
    input  wire [5-1:0]              S_AXI_MCU_DMA_AWID,
    input  wire [              31:0] S_AXI_MCU_DMA_AWADDR,
    input  wire [               2:0] S_AXI_MCU_DMA_AWSIZE,
    input  wire [               2:0] S_AXI_MCU_DMA_AWPROT,
    input  wire [               7:0] S_AXI_MCU_DMA_AWLEN,
    input  wire [               1:0] S_AXI_MCU_DMA_AWBURST,


    input  wire                      S_AXI_MCU_DMA_WVALID,
    output wire                      S_AXI_MCU_DMA_WREADY,
    input  wire [63:0]               S_AXI_MCU_DMA_WDATA,
    input  wire [ 7:0]               S_AXI_MCU_DMA_WSTRB,
    input  wire                      S_AXI_MCU_DMA_WLAST,

    output wire                      S_AXI_MCU_DMA_BVALID,
    input  wire                      S_AXI_MCU_DMA_BREADY,
    output wire [               1:0] S_AXI_MCU_DMA_BRESP,
    output wire [5-1:0]              S_AXI_MCU_DMA_BID,

    // AXI Read CHANNELS
    input  wire                      S_AXI_MCU_DMA_ARVALID,
    output wire                      S_AXI_MCU_DMA_ARREADY,
    input  wire [5-1:0]              S_AXI_MCU_DMA_ARID,
    input  wire [              31:0] S_AXI_MCU_DMA_ARADDR,
    input  wire [               2:0] S_AXI_MCU_DMA_ARSIZE,
    input  wire [               2:0] S_AXI_MCU_DMA_ARPROT,
    input  wire [               7:0] S_AXI_MCU_DMA_ARLEN,
    input  wire [               1:0] S_AXI_MCU_DMA_ARBURST,

    output wire                      S_AXI_MCU_DMA_RVALID,
    input  wire                      S_AXI_MCU_DMA_RREADY,
    output wire [5-1:0]              S_AXI_MCU_DMA_RID,
    output wire [              63:0] S_AXI_MCU_DMA_RDATA,
    output wire [               1:0] S_AXI_MCU_DMA_RRESP,
    output wire                      S_AXI_MCU_DMA_RLAST
    );

caliptra_ss_top_fpga ss_wrapper (
    
    .core_clk(core_clk),
    // Caliptra AXI Interface
    .S_AXI_CALIPTRA_AWADDR(S_AXI_CALIPTRA_AWADDR),
    .S_AXI_CALIPTRA_AWBURST(S_AXI_CALIPTRA_AWBURST),
    .S_AXI_CALIPTRA_AWSIZE(S_AXI_CALIPTRA_AWSIZE),
    .S_AXI_CALIPTRA_AWLEN(S_AXI_CALIPTRA_AWLEN),
    .S_AXI_CALIPTRA_AWUSER(S_AXI_CALIPTRA_AWUSER),
    .S_AXI_CALIPTRA_AWID(S_AXI_CALIPTRA_AWID),
    .S_AXI_CALIPTRA_AWLOCK(S_AXI_CALIPTRA_AWLOCK),
    .S_AXI_CALIPTRA_AWVALID(S_AXI_CALIPTRA_AWVALID),
    .S_AXI_CALIPTRA_AWREADY(S_AXI_CALIPTRA_AWREADY),
    // W
    .S_AXI_CALIPTRA_WDATA(S_AXI_CALIPTRA_WDATA),
    .S_AXI_CALIPTRA_WSTRB(S_AXI_CALIPTRA_WSTRB),
    .S_AXI_CALIPTRA_WVALID(S_AXI_CALIPTRA_WVALID),
    .S_AXI_CALIPTRA_WREADY(S_AXI_CALIPTRA_WREADY),
    .S_AXI_CALIPTRA_WLAST(S_AXI_CALIPTRA_WLAST),
    // B
    .S_AXI_CALIPTRA_BRESP(S_AXI_CALIPTRA_BRESP),
    .S_AXI_CALIPTRA_BID(S_AXI_CALIPTRA_BID),
    .S_AXI_CALIPTRA_BVALID(S_AXI_CALIPTRA_BVALID),
    .S_AXI_CALIPTRA_BREADY(S_AXI_CALIPTRA_BREADY),
    // AR
    .S_AXI_CALIPTRA_ARADDR(S_AXI_CALIPTRA_ARADDR),
    .S_AXI_CALIPTRA_ARBURST(S_AXI_CALIPTRA_ARBURST),
    .S_AXI_CALIPTRA_ARSIZE(S_AXI_CALIPTRA_ARSIZE),
    .S_AXI_CALIPTRA_ARLEN(S_AXI_CALIPTRA_ARLEN),
    .S_AXI_CALIPTRA_ARUSER(S_AXI_CALIPTRA_ARUSER),
    .S_AXI_CALIPTRA_ARID(S_AXI_CALIPTRA_ARID),
    .S_AXI_CALIPTRA_ARLOCK(S_AXI_CALIPTRA_ARLOCK),
    .S_AXI_CALIPTRA_ARVALID(S_AXI_CALIPTRA_ARVALID),
    .S_AXI_CALIPTRA_ARREADY(S_AXI_CALIPTRA_ARREADY),
    // R
    .S_AXI_CALIPTRA_RDATA(S_AXI_CALIPTRA_RDATA),
    .S_AXI_CALIPTRA_RRESP(S_AXI_CALIPTRA_RRESP),
    .S_AXI_CALIPTRA_RID(S_AXI_CALIPTRA_RID),
    .S_AXI_CALIPTRA_RLAST(S_AXI_CALIPTRA_RLAST),
    .S_AXI_CALIPTRA_RVALID(S_AXI_CALIPTRA_RVALID),
    .S_AXI_CALIPTRA_RREADY(S_AXI_CALIPTRA_RREADY),

    //-------------------------- LSU AXI signals--------------------------
    // AXI Write Channels
    .M_AXI_MCU_LSU_AWVALID(M_AXI_MCU_LSU_AWVALID),
    .M_AXI_MCU_LSU_AWREADY(M_AXI_MCU_LSU_AWREADY),
    .M_AXI_MCU_LSU_AWID(M_AXI_MCU_LSU_AWID),
    .M_AXI_MCU_LSU_AWADDR(M_AXI_MCU_LSU_AWADDR),
    .M_AXI_MCU_LSU_AWREGION(M_AXI_MCU_LSU_AWREGION),
    .M_AXI_MCU_LSU_AWLEN(M_AXI_MCU_LSU_AWLEN),
    .M_AXI_MCU_LSU_AWSIZE(M_AXI_MCU_LSU_AWSIZE),
    .M_AXI_MCU_LSU_AWBURST(M_AXI_MCU_LSU_AWBURST),
    .M_AXI_MCU_LSU_AWLOCK(M_AXI_MCU_LSU_AWLOCK),
    .M_AXI_MCU_LSU_AWCACHE(M_AXI_MCU_LSU_AWCACHE),
    .M_AXI_MCU_LSU_AWPROT(M_AXI_MCU_LSU_AWPROT),
    .M_AXI_MCU_LSU_AWQOS(M_AXI_MCU_LSU_AWQOS),

    .M_AXI_MCU_LSU_WVALID(M_AXI_MCU_LSU_WVALID),
    .M_AXI_MCU_LSU_WREADY(M_AXI_MCU_LSU_WREADY),
    .M_AXI_MCU_LSU_WDATA(M_AXI_MCU_LSU_WDATA),
    .M_AXI_MCU_LSU_WSTRB(M_AXI_MCU_LSU_WSTRB),
    .M_AXI_MCU_LSU_WLAST(M_AXI_MCU_LSU_WLAST),

    .M_AXI_MCU_LSU_BVALID(M_AXI_MCU_LSU_BVALID),
    .M_AXI_MCU_LSU_BREADY(M_AXI_MCU_LSU_BREADY),
    .M_AXI_MCU_LSU_BRESP(M_AXI_MCU_LSU_BRESP),
    .M_AXI_MCU_LSU_BID(M_AXI_MCU_LSU_BID),

    // AXI Read Channels
    .M_AXI_MCU_LSU_ARVALID(M_AXI_MCU_LSU_ARVALID),
    .M_AXI_MCU_LSU_ARREADY(M_AXI_MCU_LSU_ARREADY),
    .M_AXI_MCU_LSU_ARID(M_AXI_MCU_LSU_ARID),
    .M_AXI_MCU_LSU_ARADDR(M_AXI_MCU_LSU_ARADDR),
    .M_AXI_MCU_LSU_ARREGION(M_AXI_MCU_LSU_ARREGION),
    .M_AXI_MCU_LSU_ARLEN(M_AXI_MCU_LSU_ARLEN),
    .M_AXI_MCU_LSU_ARSIZE(M_AXI_MCU_LSU_ARSIZE),
    .M_AXI_MCU_LSU_ARBURST(M_AXI_MCU_LSU_ARBURST),
    .M_AXI_MCU_LSU_ARLOCK(M_AXI_MCU_LSU_ARLOCK),
    .M_AXI_MCU_LSU_ARCACHE(M_AXI_MCU_LSU_ARCACHE),
    .M_AXI_MCU_LSU_ARPROT(M_AXI_MCU_LSU_ARPROT),
    .M_AXI_MCU_LSU_ARQOS(M_AXI_MCU_LSU_ARQOS),

    .M_AXI_MCU_LSU_RVALID(M_AXI_MCU_LSU_RVALID),
    .M_AXI_MCU_LSU_RREADY(M_AXI_MCU_LSU_RREADY),
    .M_AXI_MCU_LSU_RID(M_AXI_MCU_LSU_RID),
    .M_AXI_MCU_LSU_RDATA(M_AXI_MCU_LSU_RDATA),
    .M_AXI_MCU_LSU_RRESP(M_AXI_MCU_LSU_RRESP),
    .M_AXI_MCU_LSU_RLAST(M_AXI_MCU_LSU_RLAST),

    //-------------------------- IFU AXI signals--------------------------
    // AXI Write Channels
    .M_AXI_MCU_IFU_AWVALID(M_AXI_MCU_IFU_AWVALID),
    .M_AXI_MCU_IFU_AWREADY(M_AXI_MCU_IFU_AWREADY),
    .M_AXI_MCU_IFU_AWID(M_AXI_MCU_IFU_AWID),
    .M_AXI_MCU_IFU_AWADDR(M_AXI_MCU_IFU_AWADDR),
    .M_AXI_MCU_IFU_AWREGION(M_AXI_MCU_IFU_AWREGION),
    .M_AXI_MCU_IFU_AWLEN(M_AXI_MCU_IFU_AWLEN),
    .M_AXI_MCU_IFU_AWSIZE(M_AXI_MCU_IFU_AWSIZE),
    .M_AXI_MCU_IFU_AWBURST(M_AXI_MCU_IFU_AWBURST),
    .M_AXI_MCU_IFU_AWLOCK(M_AXI_MCU_IFU_AWLOCK),
    .M_AXI_MCU_IFU_AWCACHE(M_AXI_MCU_IFU_AWCACHE),
    .M_AXI_MCU_IFU_AWPROT(M_AXI_MCU_IFU_AWPROT),
    .M_AXI_MCU_IFU_AWQOS(M_AXI_MCU_IFU_AWQOS),

    .M_AXI_MCU_IFU_WVALID(M_AXI_MCU_IFU_WVALID),
    .M_AXI_MCU_IFU_WREADY(M_AXI_MCU_IFU_WREADY),
    .M_AXI_MCU_IFU_WDATA(M_AXI_MCU_IFU_WDATA),
    .M_AXI_MCU_IFU_WSTRB(M_AXI_MCU_IFU_WSTRB),
    .M_AXI_MCU_IFU_WLAST(M_AXI_MCU_IFU_WLAST),

    .M_AXI_MCU_IFU_BVALID(M_AXI_MCU_IFU_BVALID),
    .M_AXI_MCU_IFU_BREADY(M_AXI_MCU_IFU_BREADY),
    .M_AXI_MCU_IFU_BRESP(M_AXI_MCU_IFU_BRESP),
    .M_AXI_MCU_IFU_BID(M_AXI_MCU_IFU_BID),

    // AXI Read Channels
    .M_AXI_MCU_IFU_ARVALID(M_AXI_MCU_IFU_ARVALID),
    .M_AXI_MCU_IFU_ARREADY(M_AXI_MCU_IFU_ARREADY),
    .M_AXI_MCU_IFU_ARID(M_AXI_MCU_IFU_ARID),
    .M_AXI_MCU_IFU_ARADDR(M_AXI_MCU_IFU_ARADDR),
    .M_AXI_MCU_IFU_ARREGION(M_AXI_MCU_IFU_ARREGION),
    .M_AXI_MCU_IFU_ARLEN(M_AXI_MCU_IFU_ARLEN),
    .M_AXI_MCU_IFU_ARSIZE(M_AXI_MCU_IFU_ARSIZE),
    .M_AXI_MCU_IFU_ARBURST(M_AXI_MCU_IFU_ARBURST),
    .M_AXI_MCU_IFU_ARLOCK(M_AXI_MCU_IFU_ARLOCK),
    .M_AXI_MCU_IFU_ARCACHE(M_AXI_MCU_IFU_ARCACHE),
    .M_AXI_MCU_IFU_ARPROT(M_AXI_MCU_IFU_ARPROT),
    .M_AXI_MCU_IFU_ARQOS(M_AXI_MCU_IFU_ARQOS),

    .M_AXI_MCU_IFU_RVALID(M_AXI_MCU_IFU_RVALID),
    .M_AXI_MCU_IFU_RREADY(M_AXI_MCU_IFU_RREADY),
    .M_AXI_MCU_IFU_RID(M_AXI_MCU_IFU_RID),
    .M_AXI_MCU_IFU_RDATA(M_AXI_MCU_IFU_RDATA),
    .M_AXI_MCU_IFU_RRESP(M_AXI_MCU_IFU_RRESP),
    .M_AXI_MCU_IFU_RLAST(M_AXI_MCU_IFU_RLAST),

    //-------------------------- SB AXI signals--------------------------
    // AXI Write Channels
    .sb_axi_awvalid(sb_axi_awvalid),
    .sb_axi_awready(sb_axi_awready),
    .sb_axi_awid(sb_axi_awid),
    .sb_axi_awaddr(sb_axi_awaddr),
    .sb_axi_awregion(sb_axi_awregion),
    .sb_axi_awlen(sb_axi_awlen),
    .sb_axi_awsize(sb_axi_awsize),
    .sb_axi_awburst(sb_axi_awburst),
    .sb_axi_awlock(sb_axi_awlock),
    .sb_axi_awcache(sb_axi_awcache),
    .sb_axi_awprot(sb_axi_awprot),
    .sb_axi_awqos(sb_axi_awqos),

    .sb_axi_wvalid(sb_axi_wvalid),
    .sb_axi_wready(sb_axi_wready),
    .sb_axi_wdata(sb_axi_wdata),
    .sb_axi_wstrb(sb_axi_wstrb),
    .sb_axi_wlast(sb_axi_wlast),

    .sb_axi_bvalid(sb_axi_bvalid),
    .sb_axi_bready(sb_axi_bready),
    .sb_axi_bresp(sb_axi_bresp),
    .sb_axi_bid(sb_axi_bid),

    // AXI Read Channels
    .sb_axi_arvalid(sb_axi_arvalid),
    .sb_axi_arready(sb_axi_arready),
    .sb_axi_arid(sb_axi_arid),
    .sb_axi_araddr(sb_axi_araddr),
    .sb_axi_arregion(sb_axi_arregion),
    .sb_axi_arlen(sb_axi_arlen),
    .sb_axi_arsize(sb_axi_arsize),
    .sb_axi_arburst(sb_axi_arburst),
    .sb_axi_arlock(sb_axi_arlock),
    .sb_axi_arcache(sb_axi_arcache),
    .sb_axi_arprot(sb_axi_arprot),
    .sb_axi_arqos(sb_axi_arqos),

    .sb_axi_rvalid(sb_axi_rvalid),
    .sb_axi_rready(sb_axi_rready),
    .sb_axi_rid(sb_axi_rid),
    .sb_axi_rdata(sb_axi_rdata),
    .sb_axi_rresp(sb_axi_rresp),
    .sb_axi_rlast(sb_axi_rlast),

    //-------------------------- DMA AXI signals--------------------------
    // AXI Write Channels
    .S_AXI_MCU_DMA_AWVALID(S_AXI_MCU_DMA_AWVALID),
    .S_AXI_MCU_DMA_AWREADY(S_AXI_MCU_DMA_AWREADY),
    .S_AXI_MCU_DMA_AWID(S_AXI_MCU_DMA_AWID),
    .S_AXI_MCU_DMA_AWADDR(S_AXI_MCU_DMA_AWADDR),
    .S_AXI_MCU_DMA_AWSIZE(S_AXI_MCU_DMA_AWSIZE),
    .S_AXI_MCU_DMA_AWPROT(S_AXI_MCU_DMA_AWPROT),
    .S_AXI_MCU_DMA_AWLEN(S_AXI_MCU_DMA_AWLEN),
    .S_AXI_MCU_DMA_AWBURST(S_AXI_MCU_DMA_AWBURST),


    .S_AXI_MCU_DMA_WVALID(S_AXI_MCU_DMA_WVALID),
    .S_AXI_MCU_DMA_WREADY(S_AXI_MCU_DMA_WREADY),
    .S_AXI_MCU_DMA_WDATA(S_AXI_MCU_DMA_WDATA),
    .S_AXI_MCU_DMA_WSTRB(S_AXI_MCU_DMA_WSTRB),
    .S_AXI_MCU_DMA_WLAST(S_AXI_MCU_DMA_WLAST),

    .S_AXI_MCU_DMA_BVALID(S_AXI_MCU_DMA_BVALID),
    .S_AXI_MCU_DMA_BREADY(S_AXI_MCU_DMA_BREADY),
    .S_AXI_MCU_DMA_BRESP(S_AXI_MCU_DMA_BRESP),
    .S_AXI_MCU_DMA_BID(S_AXI_MCU_DMA_BID),

    // AXI Read CHANNELS
    .S_AXI_MCU_DMA_ARVALID(S_AXI_MCU_DMA_ARVALID),
    .S_AXI_MCU_DMA_ARREADY(S_AXI_MCU_DMA_ARREADY),
    .S_AXI_MCU_DMA_ARID(S_AXI_MCU_DMA_ARID),
    .S_AXI_MCU_DMA_ARADDR(S_AXI_MCU_DMA_ARADDR),
    .S_AXI_MCU_DMA_ARSIZE(S_AXI_MCU_DMA_ARSIZE),
    .S_AXI_MCU_DMA_ARPROT(S_AXI_MCU_DMA_ARPROT),
    .S_AXI_MCU_DMA_ARLEN(S_AXI_MCU_DMA_ARLEN),
    .S_AXI_MCU_DMA_ARBURST(S_AXI_MCU_DMA_ARBURST),

    .S_AXI_MCU_DMA_RVALID(S_AXI_MCU_DMA_RVALID),
    .S_AXI_MCU_DMA_RREADY(S_AXI_MCU_DMA_RREADY),
    .S_AXI_MCU_DMA_RID(S_AXI_MCU_DMA_RID),
    .S_AXI_MCU_DMA_RDATA(S_AXI_MCU_DMA_RDATA),
    .S_AXI_MCU_DMA_RRESP(S_AXI_MCU_DMA_RRESP),
    .S_AXI_MCU_DMA_RLAST(S_AXI_MCU_DMA_RLAST)
);

endmodule