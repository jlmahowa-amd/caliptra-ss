//********************************************************************************
// SPDX-License-Identifier: Apache-2.0
// Copyright (c) 2023 Antmicro <www.antmicro.com>
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//********************************************************************************

module mcu_top
    import mcu_el2_pkg::*;
#(
    `include "mcu_el2_param.vh"
) (
    input logic        clk,
    input logic        rst_l,
    input logic        dbg_rst_l,
    input logic [31:1] rst_vec,
    input logic        nmi_int,
    input logic [31:1] nmi_vec,
    input logic [31:1] jtag_id,


    output logic [31:0] trace_rv_i_insn_ip,
    output logic [31:0] trace_rv_i_address_ip,
    output logic        trace_rv_i_valid_ip,
    output logic        trace_rv_i_exception_ip,
    output logic [ 4:0] trace_rv_i_ecause_ip,
    output logic        trace_rv_i_interrupt_ip,
    output logic [31:0] trace_rv_i_tval_ip,

    // Bus signals
`ifdef MCU_RV_BUILD_AXI4
    //-------------------------- LSU AXI signals--------------------------
    // AXI Write Channels
    output logic                      lsu_axi_awvalid,
    input  logic                      lsu_axi_awready,
    output logic [mcu_pt.LSU_BUS_TAG-1:0] lsu_axi_awid,
    output logic [              31:0] lsu_axi_awaddr,
    output logic [               3:0] lsu_axi_awregion,
    output logic [               7:0] lsu_axi_awlen,
    output logic [               2:0] lsu_axi_awsize,
    output logic [               1:0] lsu_axi_awburst,
    output logic                      lsu_axi_awlock,
    output logic [               3:0] lsu_axi_awcache,
    output logic [               2:0] lsu_axi_awprot,
    output logic [               3:0] lsu_axi_awqos,

    output logic        lsu_axi_wvalid,
    input  logic        lsu_axi_wready,
    output logic [63:0] lsu_axi_wdata,
    output logic [ 7:0] lsu_axi_wstrb,
    output logic        lsu_axi_wlast,

    input  logic                      lsu_axi_bvalid,
    output logic                      lsu_axi_bready,
    input  logic [               1:0] lsu_axi_bresp,
    input  logic [mcu_pt.LSU_BUS_TAG-1:0] lsu_axi_bid,

    // AXI Read Channels
    output logic                      lsu_axi_arvalid,
    input  logic                      lsu_axi_arready,
    output logic [mcu_pt.LSU_BUS_TAG-1:0] lsu_axi_arid,
    output logic [              31:0] lsu_axi_araddr,
    output logic [               3:0] lsu_axi_arregion,
    output logic [               7:0] lsu_axi_arlen,
    output logic [               2:0] lsu_axi_arsize,
    output logic [               1:0] lsu_axi_arburst,
    output logic                      lsu_axi_arlock,
    output logic [               3:0] lsu_axi_arcache,
    output logic [               2:0] lsu_axi_arprot,
    output logic [               3:0] lsu_axi_arqos,

    input  logic                      lsu_axi_rvalid,
    output logic                      lsu_axi_rready,
    input  logic [mcu_pt.LSU_BUS_TAG-1:0] lsu_axi_rid,
    input  logic [              63:0] lsu_axi_rdata,
    input  logic [               1:0] lsu_axi_rresp,
    input  logic                      lsu_axi_rlast,

    //-------------------------- IFU AXI signals--------------------------
    // AXI Write Channels
    output logic                      ifu_axi_awvalid,
    input  logic                      ifu_axi_awready,
    output logic [mcu_pt.IFU_BUS_TAG-1:0] ifu_axi_awid,
    output logic [              31:0] ifu_axi_awaddr,
    output logic [               3:0] ifu_axi_awregion,
    output logic [               7:0] ifu_axi_awlen,
    output logic [               2:0] ifu_axi_awsize,
    output logic [               1:0] ifu_axi_awburst,
    output logic                      ifu_axi_awlock,
    output logic [               3:0] ifu_axi_awcache,
    output logic [               2:0] ifu_axi_awprot,
    output logic [               3:0] ifu_axi_awqos,

    output logic        ifu_axi_wvalid,
    input  logic        ifu_axi_wready,
    output logic [63:0] ifu_axi_wdata,
    output logic [ 7:0] ifu_axi_wstrb,
    output logic        ifu_axi_wlast,

    input  logic                      ifu_axi_bvalid,
    output logic                      ifu_axi_bready,
    input  logic [               1:0] ifu_axi_bresp,
    input  logic [mcu_pt.IFU_BUS_TAG-1:0] ifu_axi_bid,

    // AXI Read Channels
    output logic                      ifu_axi_arvalid,
    input  logic                      ifu_axi_arready,
    output logic [mcu_pt.IFU_BUS_TAG-1:0] ifu_axi_arid,
    output logic [              31:0] ifu_axi_araddr,
    output logic [               3:0] ifu_axi_arregion,
    output logic [               7:0] ifu_axi_arlen,
    output logic [               2:0] ifu_axi_arsize,
    output logic [               1:0] ifu_axi_arburst,
    output logic                      ifu_axi_arlock,
    output logic [               3:0] ifu_axi_arcache,
    output logic [               2:0] ifu_axi_arprot,
    output logic [               3:0] ifu_axi_arqos,

    input  logic                      ifu_axi_rvalid,
    output logic                      ifu_axi_rready,
    input  logic [mcu_pt.IFU_BUS_TAG-1:0] ifu_axi_rid,
    input  logic [              63:0] ifu_axi_rdata,
    input  logic [               1:0] ifu_axi_rresp,
    input  logic                      ifu_axi_rlast,

    //-------------------------- SB AXI signals--------------------------
    // AXI Write Channels
    output logic                     sb_axi_awvalid,
    input  logic                     sb_axi_awready,
    output logic [mcu_pt.SB_BUS_TAG-1:0] sb_axi_awid,
    output logic [             31:0] sb_axi_awaddr,
    output logic [              3:0] sb_axi_awregion,
    output logic [              7:0] sb_axi_awlen,
    output logic [              2:0] sb_axi_awsize,
    output logic [              1:0] sb_axi_awburst,
    output logic                     sb_axi_awlock,
    output logic [              3:0] sb_axi_awcache,
    output logic [              2:0] sb_axi_awprot,
    output logic [              3:0] sb_axi_awqos,

    output logic        sb_axi_wvalid,
    input  logic        sb_axi_wready,
    output logic [63:0] sb_axi_wdata,
    output logic [ 7:0] sb_axi_wstrb,
    output logic        sb_axi_wlast,

    input  logic                     sb_axi_bvalid,
    output logic                     sb_axi_bready,
    input  logic [              1:0] sb_axi_bresp,
    input  logic [mcu_pt.SB_BUS_TAG-1:0] sb_axi_bid,

    // AXI Read Channels
    output logic                     sb_axi_arvalid,
    input  logic                     sb_axi_arready,
    output logic [mcu_pt.SB_BUS_TAG-1:0] sb_axi_arid,
    output logic [             31:0] sb_axi_araddr,
    output logic [              3:0] sb_axi_arregion,
    output logic [              7:0] sb_axi_arlen,
    output logic [              2:0] sb_axi_arsize,
    output logic [              1:0] sb_axi_arburst,
    output logic                     sb_axi_arlock,
    output logic [              3:0] sb_axi_arcache,
    output logic [              2:0] sb_axi_arprot,
    output logic [              3:0] sb_axi_arqos,

    input  logic                     sb_axi_rvalid,
    output logic                     sb_axi_rready,
    input  logic [mcu_pt.SB_BUS_TAG-1:0] sb_axi_rid,
    input  logic [             63:0] sb_axi_rdata,
    input  logic [              1:0] sb_axi_rresp,
    input  logic                     sb_axi_rlast,

    //-------------------------- DMA AXI signals--------------------------
    // AXI Write Channels
    input  logic                      dma_axi_awvalid,
    output logic                      dma_axi_awready,
    input  logic [mcu_pt.DMA_BUS_TAG-1:0] dma_axi_awid,
    input  logic [              31:0] dma_axi_awaddr,
    input  logic [               2:0] dma_axi_awsize,
    input  logic [               2:0] dma_axi_awprot,
    input  logic [               7:0] dma_axi_awlen,
    input  logic [               1:0] dma_axi_awburst,


    input  logic        dma_axi_wvalid,
    output logic        dma_axi_wready,
    input  logic [63:0] dma_axi_wdata,
    input  logic [ 7:0] dma_axi_wstrb,
    input  logic        dma_axi_wlast,

    output logic                      dma_axi_bvalid,
    input  logic                      dma_axi_bready,
    output logic [               1:0] dma_axi_bresp,
    output logic [mcu_pt.DMA_BUS_TAG-1:0] dma_axi_bid,

    // AXI Read Channels
    input  logic                      dma_axi_arvalid,
    output logic                      dma_axi_arready,
    input  logic [mcu_pt.DMA_BUS_TAG-1:0] dma_axi_arid,
    input  logic [              31:0] dma_axi_araddr,
    input  logic [               2:0] dma_axi_arsize,
    input  logic [               2:0] dma_axi_arprot,
    input  logic [               7:0] dma_axi_arlen,
    input  logic [               1:0] dma_axi_arburst,

    output logic                      dma_axi_rvalid,
    input  logic                      dma_axi_rready,
    output logic [mcu_pt.DMA_BUS_TAG-1:0] dma_axi_rid,
    output logic [              63:0] dma_axi_rdata,
    output logic [               1:0] dma_axi_rresp,
    output logic                      dma_axi_rlast,

    //-------------------------- I3C AXI signals--------------------------
    // AXI Write Channels
    input  logic                        i3c_axi_awvalid,
    output logic                        i3c_axi_awready,
    input  logic [mcu_pt.DMA_BUS_TAG:0] i3c_axi_awid,
    input  logic [                31:0] i3c_axi_awaddr,
    input  logic [                 2:0] i3c_axi_awsize,
    input  logic [                 2:0] i3c_axi_awprot,
    input  logic [                 7:0] i3c_axi_awlen,
    input  logic [                 1:0] i3c_axi_awburst,


    input  logic        i3c_axi_wvalid,
    output logic        i3c_axi_wready,
    input  logic [63:0] i3c_axi_wdata,
    input  logic [ 7:0] i3c_axi_wstrb,
    input  logic        i3c_axi_wlast,

    output logic                        i3c_axi_bvalid,
    input  logic                        i3c_axi_bready,
    output logic [                 1:0] i3c_axi_bresp,
    output logic [mcu_pt.DMA_BUS_TAG:0] i3c_axi_bid,

    // AXI Read Channels
    input  logic                        i3c_axi_arvalid,
    output logic                        i3c_axi_arready,
    input  logic [mcu_pt.DMA_BUS_TAG:0] i3c_axi_arid,
    input  logic [                31:0] i3c_axi_araddr,
    input  logic [                 2:0] i3c_axi_arsize,
    input  logic [                 2:0] i3c_axi_arprot,
    input  logic [                 7:0] i3c_axi_arlen,
    input  logic [                 1:0] i3c_axi_arburst,

    output logic                        i3c_axi_rvalid,
    input  logic                        i3c_axi_rready,
    output logic [mcu_pt.DMA_BUS_TAG:0] i3c_axi_rid,
    output logic [                63:0] i3c_axi_rdata,
    output logic [                 1:0] i3c_axi_rresp,
    output logic                        i3c_axi_rlast,
`endif

`ifdef MCU_RV_BUILD_AHB_LITE
    //// AHB LITE BUS
    output logic [31:0] haddr,
    output logic [ 2:0] hburst,
    output logic        hmastlock,
    output logic [ 3:0] hprot,
    output logic [ 2:0] hsize,
    output logic [ 1:0] htrans,
    output logic        hwrite,

    input logic [63:0] hrdata,
    input logic        hready,
    input logic        hresp,

    // LSU AHB Master
    output logic [31:0] lsu_haddr,
    output logic [ 2:0] lsu_hburst,
    output logic        lsu_hmastlock,
    output logic [ 3:0] lsu_hprot,
    output logic [ 2:0] lsu_hsize,
    output logic [ 1:0] lsu_htrans,
    output logic        lsu_hwrite,
    output logic [63:0] lsu_hwdata,

    input  logic [63:0] lsu_hrdata,
    input  logic        lsu_hready,
    input  logic        lsu_hresp,
    // Debug Syster Bus AHB
    output logic [31:0] sb_haddr,
    output logic [ 2:0] sb_hburst,
    output logic        sb_hmastlock,
    output logic [ 3:0] sb_hprot,
    output logic [ 2:0] sb_hsize,
    output logic [ 1:0] sb_htrans,
    output logic        sb_hwrite,
    output logic [63:0] sb_hwdata,

    input logic [63:0] sb_hrdata,
    input logic        sb_hready,
    input logic        sb_hresp,

    // DMA Slave
    input logic        dma_hsel,
    input logic [31:0] dma_haddr,
    input logic [ 2:0] dma_hburst,
    input logic        dma_hmastlock,
    input logic [ 3:0] dma_hprot,
    input logic [ 2:0] dma_hsize,
    input logic [ 1:0] dma_htrans,
    input logic        dma_hwrite,
    input logic [63:0] dma_hwdata,
    input logic        dma_hreadyin,

    output logic [63:0] dma_hrdata,
    output logic        dma_hreadyout,
    output logic        dma_hresp,

    // I3C AHB bus
    input logic        i3c_hsel,
    input logic [31:0] i3c_haddr,
    input logic [ 2:0] i3c_hburst,
    input logic        i3c_hmastlock,
    input logic [ 3:0] i3c_hprot,
    input logic [ 2:0] i3c_hsize,
    input logic [ 1:0] i3c_htrans,
    input logic        i3c_hwrite,
    input logic [63:0] i3c_hwdata,
    input logic        i3c_hreadyin,

    output logic [63:0] i3c_hrdata,
    output logic        i3c_hreadyout,
    output logic        i3c_hresp,
`endif
    // clk ratio signals
    input  logic        lsu_bus_clk_en,  // Clock ratio b/w cpu core clk & AHB master interface
    input  logic        ifu_bus_clk_en,  // Clock ratio b/w cpu core clk & AHB master interface
    input  logic        dbg_bus_clk_en,  // Clock ratio b/w cpu core clk & AHB master interface
    input  logic        dma_bus_clk_en,  // Clock ratio b/w cpu core clk & AHB slave interface

    // all of these test inputs are brought to top-level; must be tied off based on usage by physical design (ie. icache or not, iccm or not, dccm or not)

    input                                   mcu_el2_ic_data_ext_in_pkt_t  [mcu_pt.ICACHE_NUM_WAYS-1:0][mcu_pt.ICACHE_BANKS_WAY-1:0] ic_data_ext_in_pkt,
    input mcu_el2_ic_tag_ext_in_pkt_t [mcu_pt.ICACHE_NUM_WAYS-1:0] ic_tag_ext_in_pkt,

    input logic                      timer_int,
    input logic                      soft_int,
    input logic [mcu_pt.PIC_TOTAL_INT:1] extintsrc_req,

    output logic dec_tlu_perfcnt0,  // toggles when slot0 perf counter 0 has an event inc
    output logic dec_tlu_perfcnt1,
    output logic dec_tlu_perfcnt2,
    output logic dec_tlu_perfcnt3,

    // ports added by the soc team
    input  logic jtag_tck,     // JTAG clk
    input  logic jtag_tms,     // JTAG TMS
    input  logic jtag_tdi,     // JTAG tdi
    input  logic jtag_trst_n,  // JTAG Reset
    output logic jtag_tdo,     // JTAG TDO
    output logic jtag_tdoEn,   // JTAG Test Data Output enable

    input logic [31:4] core_id,

    // Memory Export Interface
    output logic mem_clk,
    // ICCM
    output logic [mcu_pt.ICCM_NUM_BANKS-1:0] iccm_clken,
    output logic [mcu_pt.ICCM_NUM_BANKS-1:0] iccm_wren_bank,
    output logic [mcu_pt.ICCM_NUM_BANKS-1:0][mcu_pt.ICCM_BITS-1:mcu_pt.ICCM_BANK_INDEX_LO] iccm_addr_bank,
    output logic [mcu_pt.ICCM_NUM_BANKS-1:0][31:0] iccm_bank_wr_data,
    output logic [mcu_pt.ICCM_NUM_BANKS-1:0][mcu_pt.ICCM_ECC_WIDTH-1:0] iccm_bank_wr_ecc,
    input logic [mcu_pt.ICCM_NUM_BANKS-1:0][31:0] iccm_bank_dout,
    input logic [mcu_pt.ICCM_NUM_BANKS-1:0][mcu_pt.ICCM_ECC_WIDTH-1:0] iccm_bank_ecc,
    // DCCM
    output logic [mcu_pt.DCCM_NUM_BANKS-1:0] dccm_clken,
    output logic [mcu_pt.DCCM_NUM_BANKS-1:0] dccm_wren_bank,
    output logic [mcu_pt.DCCM_NUM_BANKS-1:0][mcu_pt.DCCM_BITS-1:(mcu_pt.DCCM_BANK_BITS+2)] dccm_addr_bank,
    output logic [mcu_pt.DCCM_NUM_BANKS-1:0][mcu_pt.DCCM_DATA_WIDTH-1:0] dccm_wr_data_bank,
    output logic [mcu_pt.DCCM_NUM_BANKS-1:0][mcu_pt.DCCM_FDATA_WIDTH-mcu_pt.DCCM_DATA_WIDTH-1:0] dccm_wr_ecc_bank,
    input logic [mcu_pt.DCCM_NUM_BANKS-1:0][mcu_pt.DCCM_DATA_WIDTH-1:0] dccm_bank_dout,
    input logic [mcu_pt.DCCM_NUM_BANKS-1:0][mcu_pt.DCCM_FDATA_WIDTH-mcu_pt.DCCM_DATA_WIDTH-1:0] dccm_bank_ecc,

    // ICCM/DCCM ECC status
    output logic iccm_ecc_single_error,
    output logic iccm_ecc_double_error,
    output logic dccm_ecc_single_error,
    output logic dccm_ecc_double_error,

    // external MPC halt/run interface
    input  logic mpc_debug_halt_req,  // Async halt request
    input  logic mpc_debug_run_req,   // Async run request
    input  logic mpc_reset_run_req,   // Run/halt after reset
    output logic mpc_debug_halt_ack,  // Halt ack
    output logic mpc_debug_run_ack,   // Run ack
    output logic debug_brkpt_status,  // debug breakpoint

    input logic i_cpu_halt_req,  // Async halt req to CPU
    output logic o_cpu_halt_ack,  // core response to halt
    output logic o_cpu_halt_status,  // 1'b1 indicates core is halted
    output logic                            o_debug_mode_status, // Core to the PMU that core is in debug mode. When core is in debug mode, the PMU should refrain from sendng a halt or run request
    input logic i_cpu_run_req,  // Async restart req to CPU
    output logic o_cpu_run_ack,  // Core response to run req
    input logic scan_mode,  // To enable scan mode
    input logic mbist_mode,  // to enable mbist

    // DMI port for uncore
    input  logic        dmi_uncore_enable,
    output logic        dmi_uncore_en,
    output logic        dmi_uncore_wr_en,
    output logic [ 6:0] dmi_uncore_addr,
    output logic [31:0] dmi_uncore_wdata,
    input  logic [31:0] dmi_uncore_rdata,

    // I3C Interface
`ifdef VERILATOR
    input  logic scl_i,
    input  logic sda_i,
    output logic scl_o,
    output logic sda_o,
    output logic sel_od_pp_o
`else
    inout  logic i3c_scl_io,
    inout  logic i3c_sda_io
`endif
);

  mcu_el2_mem_if mem_export ();
  assign mem_clk                   = mem_export.clk;
  assign dccm_clken                = mem_export.dccm_clken;
  assign dccm_wren_bank            = mem_export.dccm_wren_bank;
  assign dccm_addr_bank            = mem_export.dccm_addr_bank;
  assign dccm_wr_data_bank         = mem_export.dccm_wr_data_bank;
  assign dccm_wr_ecc_bank          = mem_export.dccm_wr_ecc_bank;
  assign mem_export.dccm_bank_dout = dccm_bank_dout;
  assign mem_export.dccm_bank_ecc  = dccm_bank_ecc;
  assign iccm_clken                = mem_export.iccm_clken;
  assign iccm_wren_bank            = mem_export.iccm_wren_bank;
  assign iccm_addr_bank            = mem_export.iccm_addr_bank;
  assign iccm_bank_wr_data         = mem_export.iccm_bank_wr_data;
  assign iccm_bank_wr_ecc          = mem_export.iccm_bank_wr_ecc;
  assign mem_export.iccm_bank_dout = iccm_bank_dout;
  assign mem_export.iccm_bank_ecc  = iccm_bank_ecc;

  mcu_el2_veer_wrapper rvtop (
      .mcu_el2_mem_export(mem_export.veer_sram_src),
      .*
  );

  i3c_wrapper #(
`ifdef MCU_RV_BUILD_AHB_LITE
    .AhbDataWidth(`CALIPTRA_AHB_HDATA_SIZE),
    .AhbAddrWidth(`CALIPTRA_SLAVE_ADDR_WIDTH(`CALIPTRA_SLAVE_SEL_I3C))
`elsif MCU_RV_BUILD_AXI4
    .AxiDataWidth(`AXI_DATA_WIDTH),
    .AxiAddrWidth(`AXI_ADDR_WIDTH),
    .AxiUserWidth(`AXI_USER_WIDTH),
    .AxiIdWidth(`AXI_ID_WIDTH)
`endif
  ) i3c (
      .clk_i(clk),
      .rst_ni(rst_l),

`ifdef MCU_RV_BUILD_AHB_LITE
      // AMBA AHB Lite Interface
      .haddr_i(i3c_haddr),
      .hburst_i(i3c_hburst),
      .hprot_i(i3c_hprot),
      .hwdata_i(i3c_hwdata),
      .hsel_i(i3c_hsel),
      .hwstrb_i(i3c_hwstrb),
      .hwrite_i(i3c_hwrite),
      .hready_i(i3c_hready),
      .htrans_i(i3c_htrans),
      .hsize_i(i3c_hsize),
      .hresp_o(i3c_hresp),
      .hreadyout_o(i3c_hreadyout),
      .hrdata_o(i3c_hrdata),
`elsif MCU_RV_BUILD_AXI4
     // AXI Read Channels
      .araddr_i(i3c_axi_araddr),
      .arburst_i(i3c_axi_arburst),
      .arsize_i(i3c_axi_arsize),
      .arlen_i(i3c_axi_arlen),
      .aruser_i(i3c_axi_aruser),
      .arid_i(i3c_axi_arid),
      .arlock_i(i3c_axi_arlock),
      .arvalid_i(i3c_axi_arvalid),
      .arready_o(i3c_axi_arready),

      .rdata_o(i3c_axi_rdata),
      .rresp_o(i3c_axi_rresp),
      .rid_o(i3c_axi_rid),
      .rlast_o(i3c_axi_rlast),
      .rvalid_o(i3c_axi_rvalid),
      .rready_i(i3c_axi_rready),

      // AXI Write Channels
      .awaddr_i(i3c_axi_awaddr),
      .awburst_i(i3c_axi_awburst),
      .awsize_i(i3c_axi_awsize),
      .awlen_i(i3c_axi_awlen),
      .awuser_i(i3c_axi_awuser),
      .awid_i(i3c_axi_awid),
      .awlock_i(i3c_axi_awlock),
      .awvalid_i(i3c_axi_awvalid),
      .awready_o(i3c_axi_awready),

      .wdata_i (i3c_axi_wdata),
      .wstrb_i (i3c_axi_wstrb),
      .wlast_i (i3c_axi_wlast),
      .wvalid_i(i3c_axi_wvalid),
      .wready_o(i3c_axi_wready),

      .bresp_o(i3c_axi_bresp),
      .bid_o(i3c_axi_bid),
      .bvalid_o(i3c_axi_bvalid),
      .bready_i(i3c_axi_bready),
`endif

`ifdef VERILATOR
      .scl_i(scl_i),
      .sda_i(sda_i),
      .scl_o(scl_o),
      .sda_o(sda_o),
      .sel_od_pp_o(sel_od_pp_o)
`else
      // I3C bus IO
      .i3c_scl_io(i3c_scl_io),
      .i3c_sda_io(i3c_sda_io)
`endif
  );

endmodule

